magic
tech sky130A
magscale 1 2
timestamp 1729097492
<< viali >>
rect 132 2309 290 2343
rect 553 2309 711 2343
rect 974 2309 1132 2343
rect 132 1289 290 1323
rect 553 1289 711 1323
rect 974 1289 1132 1323
<< metal1 >>
rect 0 2343 1264 2379
rect 0 2309 132 2343
rect 290 2309 553 2343
rect 711 2309 974 2343
rect 1132 2309 1264 2343
rect 0 2303 1264 2309
rect 0 1841 228 1847
rect 0 1781 6 1841
rect 222 1781 228 1841
rect 1110 1841 1338 1847
rect 268 1791 649 1832
rect 689 1791 1070 1832
rect 0 1775 228 1781
rect 1110 1781 1116 1841
rect 1332 1781 1338 1841
rect 1110 1775 1338 1781
rect 0 1323 1264 1329
rect 0 1289 132 1323
rect 290 1289 553 1323
rect 711 1289 974 1323
rect 1132 1289 1264 1323
rect 0 1253 1264 1289
<< via1 >>
rect 6 1781 222 1841
rect 1116 1781 1332 1841
<< metal2 >>
rect 0 1841 228 1847
rect 1110 1841 1338 1847
rect 0 1781 6 1841
rect 222 1781 1116 1841
rect 1332 1781 1338 1841
rect 0 1775 228 1781
rect 1110 1775 1338 1781
use inverter  x1 ~/ic_projects/inverter/mag
timestamp 1729092732
transform 1 0 53 0 1 1306
box -53 -53 369 1073
use inverter  x2
timestamp 1729092732
transform 1 0 474 0 1 1306
box -53 -53 369 1073
use inverter  x3
timestamp 1729092732
transform 1 0 895 0 1 1306
box -53 -53 369 1073
<< labels >>
flabel metal1 634 2361 634 2361 0 FreeSans 160 0 0 0 vdd
port 0 nsew
flabel metal1 633 1273 633 1273 0 FreeSans 160 0 0 0 gnd
port 1 nsew
flabel via1 1222 1810 1222 1810 0 FreeSans 160 0 0 0 out
port 2 nsew
<< end >>
